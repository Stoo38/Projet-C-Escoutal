library IEEE ;

library IEEE ;

library IEEE ;
