library IEEE ;
use IEEE.std_logic_1164.ALL ; --simulation d'un commentaire
use ieee.numeric_std.all; --seconde simulation
